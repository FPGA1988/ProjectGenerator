//****************************************************************************************************  
//*------------------Copyright (c) 2016 C-L-G.FPGA1988.bwang. All rights reserved---------------------
//
//                       --              It to be define                --
//                       --                    ...                      --
//                       --                    ...                      --
//                       --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : delay_module.v 
//Project Name   : gt0000
//Description    : the top module of gt0000
//Github Address : https://github.com/C-L-G/gt0000/trunk/ic/digital/rtl/gt0000_digital_top.v
//License        : CPL
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 01-07-2016 17:00(1th Fri,July,2016)
//First Author   : bwang
//Modify Date    : 02-09-2016 14:20(1th Sun,July,2016)
//Last Author    : bwang
//Version Number : 002   
//Last Commit    : 03-09-2016 14:30(1th Sun,July,2016)
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2017.06.29 - bwang - The initial version.
//*---------------------------------------------------------------------------------------------------
`timescale 1ns/1ps
module delay_module(
    //************************************************************************************************
    // 1.input and output declaration
    //************************************************************************************************
    input   wire            dly_i  ,//01   In
    output  wire            dly_o   //01   Out
);
    //************************************************************************************************
    // 2.Parameter and constant define
    //************************************************************************************************
    `define DELAY_CELL BUF_X1M_GT50
    
    parameter DELAY_LEVEL = 8   ; 
    
    
    //************************************************************************************************
    // 3.Register and wire declaration
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 3.1 the delay wire
    //------------------------------------------------------------------------------------------------   
    wire    [DELAY:00]              dly_wire    ;
    genvar                          i           ; 
    
    //------------------------------------------------------------------------------------------------
    // 3.x the test logic
    //------------------------------------------------------------------------------------------------
    //None
    
    //************************************************************************************************
    // 4.Main code
    //************************************************************************************************

    //------------------------------------------------------------------------------------------------
    // 4.1 the delay wire assignment
    //------------------------------------------------------------------------------------------------    
    assign dly_wire[0]  = dly_i;
    assign dly_o        = dly_wire[DELAY_LEVEL];

    //************************************************************************************************
    // 5.Sub module instantiation
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 5.1 the delay generate logic
    //------------------------------------------------------------------------------------------------    
    generate
        for(i=0;i<DELAY_LEVEL;i=i+1) begin : DELAY_CELL_INST
            `DELAY_CELL dly_cell_inst(.A(dly_wire[i],.Y(dly_wire[i+1]));
        end
    endgenerate

endmodule    
//****************************************************************************************************
//End of Module
//****************************************************************************************************

//****************************************************************************************************  
//*------------------Copyright (c) 2016 C-L-G.FPGA1988.bwang. All rights reserved---------------------
//
//                       --              It to be define                --
//                       --                    ...                      --
//                       --                    ...                      --
//                       --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : ecc_dec_module.v 
//Project Name   : gt0000
//Description    : the top module of gt0000
//Github Address : https://github.com/C-L-G/gt0000/trunk/ic/digital/rtl/gt0000_digital_top.v
//License        : CPL
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 01-07-2016 17:00(1th Fri,July,2016)
//First Author   : bwang
//Modify Date    : 02-09-2016 14:20(1th Sun,July,2016)
//Last Author    : bwang
//Version Number : 002   
//Last Commit    : 03-09-2016 14:30(1th Sun,July,2016)
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2017.06.29 - bwang - The initial version.
//*---------------------------------------------------------------------------------------------------
`timescale 1ns/1ps
module ecc_dec_module(
    //************************************************************************************************
    // 1.input and output declaration
    //************************************************************************************************
    input   wire    [37:00]         r   ,//the code may contain error
    output  wire    [31:00]         c    //the corrected code
);
    //************************************************************************************************
    // 2.Parameter and constant define
    //************************************************************************************************
    
    
    
    
    //************************************************************************************************
    // 3.Register and wire declaration
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 3.1 the clk wire signal
    //------------------------------------------------------------------------------------------------   
    
    
    
    //------------------------------------------------------------------------------------------------
    // 3.x the test logic
    //------------------------------------------------------------------------------------------------
    //************************************************************************************************
    // 4.Main code
    //************************************************************************************************

    //------------------------------------------------------------------------------------------------
    // 4.x the Test Logic
    //------------------------------------------------------------------------------------------------    
    //Rapid Matrix Multiplication algorithm v = v*G
    assign s[05] = r[37]^r[31]^r[30]^r[29]r[28]^r[27]^r[16]^r[15]^r[14]^r[13]^r[12]^r[11]^r[10]^r[9]^1'b0; 
    assign s[04] = r[36]^r[31]^r[26]^r[25]r[24]^r[23]^r[16]^r[15]^r[14]^r[8]^r[7]^r[6]^r[5]^r[4]^r[3]^1'b1; 
    assign s[03] = r[35]^r[30]^r[26]^r[22]r[21]^r[20]^r[13]^r[12]^r[8]^r[7]^r[6]^r[2]^r[1]^r[0]^1'b0; 
    assign s[02] = r[34]^r[29]^r[25]^r[22]r[19]^r[18]^r[16]^r[13]^r[11]^r[10]^r[8]^r[5]^r[4]^r[2]^r[1]^1'b1; 
    assign s[01] = r[33]^r[28]^r[24]^r[21]r[19]^r[17]^r[15]^r[11]^r[9]^r[7]^r[5]^r[3]^r[2]^r[0]^1'b0; 
    assign s[00] = r[32]^r[27]^r[23]^r[20]r[18]^r[17]^r[14]^r[12]^r[10]^r[9]^r[6]^r[4]^r[3]^r[1]^r[0]^1'b1; 

    assign c[37] = r[37]^( s[5] & ~s[4] & ~s[3] & ~s[2] & ~s[1] & ~s[0]);   //100000
    assign c[36] = r[36]^(~s[5] &  s[4] & ~s[3] & ~s[2] & ~s[1] & ~s[0]);   //010000
    assign c[35] = r[35]^(~s[5] & ~s[4] &  s[3] & ~s[2] & ~s[1] & ~s[0]);   //001000
    assign c[34] = r[34]^(~s[5] & ~s[4] & ~s[3] &  s[2] & ~s[1] & ~s[0]);   //000100
    assign c[33] = r[33]^(~s[5] & ~s[4] & ~s[3] & ~s[2] &  s[1] & ~s[0]);   //000010
    assign c[32] = r[32]^(~s[5] & ~s[4] & ~s[3] & ~s[2] & ~s[1] &  s[0]);   //000001
    assign c[31] = r[31]^( s[5] &  s[4] & ~s[3] & ~s[2] & ~s[1] & ~s[0]);   //110000
    assign c[30] = r[30]^( s[5] & ~s[4] &  s[3] & ~s[2] & ~s[1] & ~s[0]);   //101000
    assign c[29] = r[29]^( s[5] & ~s[4] & ~s[3] &  s[2] & ~s[1] & ~s[0]);   //100100
    assign c[28] = r[28]^( s[5] & ~s[4] & ~s[3] & ~s[2] &  s[1] & ~s[0]);   //100010
    assign c[27] = r[27]^( s[5] & ~s[4] & ~s[3] & ~s[2] & ~s[1] &  s[0]);   //100001
    assign c[26] = r[26]^(~s[5] &  s[4] &  s[3] & ~s[2] & ~s[1] & ~s[0]);   //011000
    assign c[25] = r[25]^(~s[5] &  s[4] & ~s[3] &  s[2] & ~s[1] & ~s[0]);   //010100
    assign c[24] = r[24]^(~s[5] &  s[4] & ~s[3] & ~s[2] &  s[1] & ~s[0]);   //010010
    assign c[23] = r[23]^(~s[5] &  s[4] & ~s[3] & ~s[2] & ~s[1] &  s[0]);   //010001
    assign c[22] = r[22]^(~s[5] & ~s[4] &  s[3] &  s[2] & ~s[1] & ~s[0]);   //001100
    assign c[21] = r[21]^(~s[5] & ~s[4] &  s[3] & ~s[2] &  s[1] & ~s[0]);   //001010
    assign c[20] = r[20]^(~s[5] & ~s[4] &  s[3] & ~s[2] & ~s[1] &  s[0]);   //001001
    assign c[19] = r[19]^(~s[5] & ~s[4] & ~s[3] &  s[2] &  s[1] & ~s[0]);   //000110
    assign c[18] = r[18]^(~s[5] & ~s[4] & ~s[3] &  s[2] & ~s[1] &  s[0]);   //000101
    assign c[17] = r[17]^(~s[5] & ~s[4] & ~s[3] & ~s[2] &  s[1] &  s[0]);   //0000l1
    assign c[16] = r[16]^( s[5] &  s[4] & ~s[3] &  s[2] & ~s[1] & ~s[0]);   //110100
    assign c[15] = r[15]^( s[5] &  s[4] & ~s[3] & ~s[2] &  s[1] & ~s[0]);   //110010
    assign c[14] = r[14]^( s[5] &  s[4] & ~s[3] & ~s[2] & ~s[1] &  s[0]);   //110001
    assign c[13] = r[13]^( s[5] & ~s[4] &  s[3] &  s[2] & ~s[1] & ~s[0]);   //101100
    assign c[12] = r[12]^( s[5] & ~s[4] &  s[3] & ~s[2] & ~s[1] &  s[0]);   //101001
    assign c[11] = r[11]^( s[5] & ~s[4] & ~s[3] &  s[2] &  s[1] & ~s[0]);   //100110
    assign c[10] = r[10]^( s[5] & ~s[4] & ~s[3] &  s[2] & ~s[1] &  s[0]);   //100101
    assign c[09] = r[09]^( s[5] & ~s[4] & ~s[3] & ~s[2] &  s[1] &  s[0]);   //100011
    assign c[08] = r[08]^(~s[5] &  s[4] &  s[3] &  s[2] & ~s[1] & ~s[0]);   //011100
    assign c[07] = r[07]^(~s[5] &  s[4] &  s[3] & ~s[2] &  s[1] & ~s[0]);   //011010
    assign c[06] = r[06]^(~s[5] &  s[4] &  s[3] & ~s[2] & ~s[1] &  s[0]);   //011001
    assign c[05] = r[05]^(~s[5] &  s[4] & ~s[3] &  s[2] &  s[1] & ~s[0]);   //010110
    assign c[04] = r[04]^(~s[5] &  s[4] & ~s[3] &  s[2] & ~s[1] &  s[0]);   //010101
    assign c[03] = r[03]^(~s[5] &  s[4] & ~s[3] & ~s[2] &  s[1] &  s[0]);   //010011
    assign c[02] = r[02]^(~s[5] & ~s[4] &  s[3] &  s[2] &  s[1] & ~s[0]);   //001110
    assign c[01] = r[01]^(~s[5] & ~s[4] &  s[3] &  s[2] & ~s[1] &  s[0]);   //001101
    assign c[00] = r[00]^(~s[5] & ~s[4] &  s[3] & ~s[2] &  s[1] &  s[0]);   //001011
    //************************************************************************************************
    // 5.Sub module instantiation
    //************************************************************************************************
endmodule    
//****************************************************************************************************
//End of Module
//****************************************************************************************************

//****************************************************************************************************  
//*------------------Copyright (c) 2016 C-L-G.FPGA1988.bwang. All rights reserved---------------------
//
//                       --              It to be define                --
//                       --                    ...                      --
//                       --                    ...                      --
//                       --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : gt0000_digital_top.v 
//Project Name   : gt0000
//Description    : the top module of gt0000
//Github Address : https://github.com/C-L-G/gt0000/trunk/ic/digital/rtl/gt0000_digital_top.v
//License        : CPL
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 01-07-2016 17:00(1th Fri,July,2016)
//First Author   : bwang
//Modify Date    : 02-09-2016 14:20(1th Sun,July,2016)
//Last Author    : bwang
//Version Number : 002   
//Last Commit    : 03-09-2016 14:30(1th Sun,July,2016)
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2017.06.29 - bwang - The initial version.
//*---------------------------------------------------------------------------------------------------
`timescale 1ns/1ps
module ecc_enc_module(
    input   wire    [31:00]         i   ,//the origital message
    output  wire    [37:00]         o    //the ecc code + origital data
);

    //************************************************************************************************
    // 1.input and output declaration
    //************************************************************************************************

    //************************************************************************************************
    // 2.Parameter and constant define
    //************************************************************************************************
    
    
    
    
    //************************************************************************************************
    // 3.Register and wire declaration
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 3.1 the clk wire signal
    //------------------------------------------------------------------------------------------------   
    
    
    
    //------------------------------------------------------------------------------------------------
    // 3.x the test logic
    //------------------------------------------------------------------------------------------------
    //************************************************************************************************
    // 4.Main code
    //************************************************************************************************

    //------------------------------------------------------------------------------------------------
    // 4.x the Test Logic
    //------------------------------------------------------------------------------------------------    
    //Rapid Matrix Multiplication algorithm v = v*G
    assign o[37] = i[31]^i[30]^i[29]i[28]^i[27]^i[16]^i[15]^i[14]^i[13]^i[12]^i[11]^i[10]^i[9]^1'b0; 
    assign o[36] = i[31]^i[26]^i[25]i[24]^i[23]^i[16]^i[15]^i[14]^i[8]^i[7]^i[6]^i[5]^i[4]^i[3]^1'b1; 
    assign o[35] = i[30]^i[26]^i[22]i[21]^i[20]^i[13]^i[12]^i[8]^i[7]^i[6]^i[2]^i[1]^i[0]^1'b0; 
    assign o[34] = i[29]^i[25]^i[22]i[19]^i[18]^i[16]^i[13]^i[11]^i[10]^i[8]^i[5]^i[4]^i[2]^i[1]^1'b1; 
    assign o[33] = i[28]^i[24]^i[21]i[19]^i[17]^i[15]^i[11]^i[9]^i[7]^i[5]^i[3]^i[2]^i[0]^1'b0; 
    assign o[32] = i[27]^i[23]^i[20]i[18]^i[17]^i[14]^i[12]^i[10]^i[9]^i[6]^i[4]^i[3]^i[1]^i[0]^1'b1; 
    assign o[31:0] = i[31:];
    //************************************************************************************************
    // 5.Sub module instantiation
    //************************************************************************************************
    //------------------------------------------------------------------------------------------------
    // 5.1 ecc syndrome table : G(ECC(38,32))
    //------------------------------------------------------------------------------------------------    
    /*
    000000  000000_00000000_00000000_00000000_00000000  
    100000  100000_00000000_00000000_00000000_00000000  
    010000  010000_00000000_00000000_00000000_00000000  
    001000  001000_00000000_00000000_00000000_00000000  
    000100  000100_00000000_00000000_00000000_00000000  
    000010  000010_00000000_00000000_00000000_00000000  
    000001  000001_00000000_00000000_00000000_00000000  
    110000  000000_10000000_00000000_00000000_00000000  
    101000  000000_01000000_00000000_00000000_00000000  
    100100  000000_00100000_00000000_00000000_00000000  
    100010  000000_00010000_00000000_00000000_00000000  
    100001  000000_00001000_00000000_00000000_00000000  
    011000  000000_00000100_00000000_00000000_00000000  
    010100  000000_00000010_00000000_00000000_00000000  
    010010  000000_00000001_00000000_00000000_00000000  
    010001  000000_00000000_10000000_00000000_00000000  
    001100  000000_00000000_01000000_00000000_00000000  
    001010  000000_00000000_00100000_00000000_00000000  
    001001  000000_00000000_00010000_00000000_00000000  
    000110  000000_00000000_00001000_00000000_00000000  
    000101  000000_00000000_00000100_00000000_00000000  
    000011  000000_00000000_00000010_00000000_00000000  
    110100  000000_00000000_00000001_00000000_00000000  
    110010  000000_00000000_00000000_10000000_00000000  
    110001  000000_00000000_00000000_01000000_00000000  
    101100  000000_00000000_00000000_00100000_00000000  
    101001  000000_00000000_00000000_00010000_00000000  
    100110  000000_00000000_00000000_00001000_00000000  
    100101  000000_00000000_00000000_00000100_00000000  
    100011  000000_00000000_00000000_00000010_00000000  
    011100  000000_00000000_00000000_00000001_00000000  
    011010  000000_00000000_00000000_00000000_10000000  
    011001  000000_00000000_00000000_00000000_01000000  
    011001  000000_00000000_00000000_00000000_01000000  
    010110  000000_00000000_00000000_00000000_00100000  
    010101  000000_00000000_00000000_00000000_00010000  
    010011  000000_00000000_00000000_00000000_00001000  
    001110  000000_00000000_00000000_00000000_00000100  
    001101  000000_00000000_00000000_00000000_00000010  
    001011  000000_00000000_00000000_00000000_00000001  
    101010  000000_00000000_00000000_00000000_0000000010 virtual 
    111111  000000_00000000_00000000_00000000_0000000001 virtual 
    */
endmodule    
//****************************************************************************************************
//End of Module
//****************************************************************************************************


//****************************************************************************************************  
//*------------------Copyright (c) 2016 C-L-G.FPGA1988.bwang. All rights reserved---------------------
//
//                   --              It to be define                --
//                   --                    ...                      --
//                   --                    ...                      --
//                   --                    ...                      --
//**************************************************************************************************** 
//File Information
//**************************************************************************************************** 
//File Name      : digital_top.v 
//Project Name   : gt0000
//Description    : the top module of gt0000
//Github Address : https://github.com/C-L-G/gt0000/trunk/ic/digital/rtl/digital_top.v
//License        : CPL
//**************************************************************************************************** 
//Version Information
//**************************************************************************************************** 
//Create Date    : 2017.07.18
//First Author   : bwang
//Modify Date    : 2017.07.18
//Last Author    : bwang
//Version Number : 002   
//Last Commit    : 2017.07.18
//**************************************************************************************************** 
//Change History(latest change first)
//yyyy.mm.dd - Author - Your log of change
//**************************************************************************************************** 
//2017.07.18 - bwang - Add the clock switch test logic,rename the clk gen module to clk gen top.
//2017.07.18 - bwang - Add the system auxiliary module,add the test logic.
//2017.07.18 - bwang - The initial version.
//*---------------------------------------------------------------------------------------------------

